module UART_RX(CLK50MHz, DATA);
	input CLK50MHz;
	output [7:0] DATA;
	
	
	
endmodule
