
module niosSystem (
	clk_clk,
	reset_reset_n,
	green_leds_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	green_leds_export;
endmodule
